module iramHRM(CLK, RESET, ADDR, Q);
  input           CLK;
  input           RESET;
  input  [9:0]  ADDR; // Enlargened for PC
  output [15:0] Q;

  reg     [15:0] mem[0:511]; // instruction memory with 16 bit entries

  wire    [8:0]  saddr;
  integer        i;


  assign saddr = ADDR[9:1];
  assign Q = mem[saddr];

  always @(posedge CLK) begin
     if(RESET) begin
        mem[0]   <= 16'b1111000000000001;    // SUB R0, R0, R0
        mem[1]   <= 16'b1111000000001000;    // ADD R1, R0, R0
        mem[2]   <= 16'b1111000000010000;    // ADD R2, R0, R0
        mem[3]   <= 16'b1111000000011000;    // ADD R3, R0, R0
        mem[4]   <= 16'b0100000000110111;    // SB R0, -9(R0)
        mem[5]   <= 16'b0010000100110110;    // LB R4, -10(R0)
        mem[6]   <= 16'b1001000100000001;    // BNE R4, R0, continue_mini_if[1]
        mem[7]   <= 16'b0001000000000100;    // JUMP while[4]
        mem[8]   <= 16'b1111001000111100;    // SLL R7, R1
        mem[9]   <= 16'b1111111000111100;    // SLL R7, R7
        mem[10]  <= 16'b1111111000111100;    // SLL R7, R7
        mem[11]  <= 16'b1111111000111100;    // SLL R7, R7
        mem[12]  <= 16'b1111111010111000;    // ADD R7, R7, R2
        mem[13]  <= 16'b0101111111011110;    // ADDI R7, R7, 30
        mem[14]  <= 16'b0101111111011110;    // ADDI R7, R7, 30
        mem[15]  <= 16'b0101111111000100;    // ADDI R7, R7, 4
        mem[16]  <= 16'b0010111101000000;    // LB R5, 0(R7)
        mem[17]  <= 16'b0101000110111111;    // ADDI R6, R0, -1
        mem[18]  <= 16'b1111110000110011;    // SRL R6, R6
        mem[19]  <= 16'b1111101110101101;    // AND R5, R5, R6
        mem[20]  <= 16'b0100111101000000;    // SB R5, 0(R7)
        mem[21]  <= 16'b0101000111000111;    // ADDI R7, R0, 7
        mem[22]  <= 16'b1001111100000100;    // BNE R4, R7, elif_1[4]
        mem[23]  <= 16'b0101010111111111;    // ADDI R7, R2, -1
        mem[24]  <= 16'b1011111000000010;    // BLTZ R7, elif_1[2]
        mem[25]  <= 16'b0101010010111111;    // ADDI R2, R2, -1
        mem[26]  <= 16'b0001000001011000;    // JUMP elif_done[88]
        mem[27]  <= 16'b0101000111000101;    // ADDI R7, R0, 5
        mem[28]  <= 16'b1001111100000100;    // BNE R4, R7, elif_2[4]
        mem[29]  <= 16'b0101010111110001;    // ADDI R7, R2, -15
        mem[30]  <= 16'b1010111000000010;    // BGEZ R7, elif_2[2]
        mem[31]  <= 16'b0101010010000001;    // ADDI R2, R2, 1
        mem[32]  <= 16'b0001000001011000;    // JUMP elif_done[88]
        mem[33]  <= 16'b0101000111000100;    // ADDI R7, R0, 4
        mem[34]  <= 16'b1001111100000100;    // BNE R4, R7, elif_3[4]
        mem[35]  <= 16'b0101001111111111;    // ADDI R7, R1, -1
        mem[36]  <= 16'b1011111000000010;    // BLTZ R7, elif_3[2]
        mem[37]  <= 16'b0101001001111111;    // ADDI R1, R1, -1
        mem[38]  <= 16'b0001000001011000;    // JUMP elif_done[88]
        mem[39]  <= 16'b0101000111000110;    // ADDI R7, R0, 6
        mem[40]  <= 16'b1001111100000100;    // BNE R4, R7, elif_4[4]
        mem[41]  <= 16'b0101001111111101;    // ADDI R7, R1, -3
        mem[42]  <= 16'b1010111000000010;    // BGEZ R7, elif_4[2]
        mem[43]  <= 16'b0101001001000001;    // ADDI R1, R1, 1
        mem[44]  <= 16'b0001000001011000;    // JUMP elif_done[88]
        mem[45]  <= 16'b0101000111000001;    // ADDI R7, R0, 1
        mem[46]  <= 16'b1000111100000001;    // BEQ R4, R7, continue_elif_4[1]
        mem[47]  <= 16'b0001000001001100;    // JUMP elif_5[76]
        mem[48]  <= 16'b1111001000111100;    // SLL R7, R1
        mem[49]  <= 16'b1111111000111100;    // SLL R7, R7
        mem[50]  <= 16'b1111111000111100;    // SLL R7, R7
        mem[51]  <= 16'b1111111000111100;    // SLL R7, R7
        mem[52]  <= 16'b1111111010111000;    // ADD R7, R7, R2
        mem[53]  <= 16'b0101111111011110;    // ADDI R7, R7, 30
        mem[54]  <= 16'b0101111111011110;    // ADDI R7, R7, 30
        mem[55]  <= 16'b0101111111000100;    // ADDI R7, R7, 4
        mem[56]  <= 16'b0010111110000000;    // LB R6, 0(R7)
        mem[57]  <= 16'b1111110000110100;    // SLL R6, R6
        mem[58]  <= 16'b1111110000110011;    // SRL R6, R6
        mem[59]  <= 16'b0101110110100010;    // ADDI R6, R6, -30
        mem[60]  <= 16'b0101110110100010;    // ADDI R6, R6, -30
        mem[61]  <= 16'b0101110110111101;    // ADDI R6, R6, -3
        mem[62]  <= 16'b1001000110000100;    // BNE R6, R0, not_question[4]
        mem[63]  <= 16'b0101000110010000;    // ADDI R6, R0, 16
        mem[64]  <= 16'b0101110110010000;    // ADDI R6, R6, 16
        mem[65]  <= 16'b0100111110000000;    // SB R6, 0(R7)
        mem[66]  <= 16'b0001000001011000;    // JUMP elif_done[88]
        mem[67]  <= 16'b0010111110000000;    // LB R6, 0(R7)
        mem[68]  <= 16'b0101110110110000;    // ADDI R6, R6, -16
        mem[69]  <= 16'b0101110110110000;    // ADDI R6, R6, -16
        mem[70]  <= 16'b1001000110000101;    // BNE R6, R0, elif_5[5]
        mem[71]  <= 16'b0101000110011110;    // ADDI R6, R0, 30
        mem[72]  <= 16'b0101110110011110;    // ADDI R6, R6, 30
        mem[73]  <= 16'b0101110110000011;    // ADDI R6, R6, 3
        mem[74]  <= 16'b0100111110000000;    // SB R6, 0(R7)
        mem[75]  <= 16'b0001000001011000;    // JUMP elif_done[88]
        mem[76]  <= 16'b0101000111000010;    // ADDI R7, R0, 2
        mem[77]  <= 16'b1001111100001010;    // BNE R4, R7, elif_done[10]
        mem[78]  <= 16'b1111001000111100;    // SLL R7, R1
        mem[79]  <= 16'b1111111000111100;    // SLL R7, R7
        mem[80]  <= 16'b1111111000111100;    // SLL R7, R7
        mem[81]  <= 16'b1111111000111100;    // SLL R7, R7
        mem[82]  <= 16'b1111111010111000;    // ADD R7, R7, R2
        mem[83]  <= 16'b0010111110000000;    // LB R6, 0(R7)
        mem[84]  <= 16'b0101111111011110;    // ADDI R7, R7, 30
        mem[85]  <= 16'b0101111111011110;    // ADDI R7, R7, 30
        mem[86]  <= 16'b0101111111000100;    // ADDI R7, R7, 4
        mem[87]  <= 16'b0100111110000000;    // SB R6, 0(R7)
        mem[88]  <= 16'b1111001000111100;    // SLL R7, R1
        mem[89]  <= 16'b1111111000111100;    // SLL R7, R7
        mem[90]  <= 16'b1111111000111100;    // SLL R7, R7
        mem[91]  <= 16'b1111111000111100;    // SLL R7, R7
        mem[92]  <= 16'b1111111010111000;    // ADD R7, R7, R2
        mem[93]  <= 16'b0101111111011110;    // ADDI R7, R7, 30
        mem[94]  <= 16'b0101111111011110;    // ADDI R7, R7, 30
        mem[95]  <= 16'b0101111111000100;    // ADDI R7, R7, 4
        mem[96]  <= 16'b0010111110000000;    // LB R6, 0(R7)
        mem[97]  <= 16'b0111110110111111;    // ORI R6, R6, -1
        mem[98]  <= 16'b0100111110000000;    // SB R6, 0(R7)
        mem[99]  <= 16'b0101000110001111;    // ADDI R6, R0, 15
        mem[100] <= 16'b0100000110110111;    // SB R6, -9(R0)
        mem[101] <= 16'b0001000000000100;    // JUMP while[4]

       for(i = 102; i < 512; i = i + 1) begin // Updated PC limit
          mem[i] <= 16'b0000000000000000;
        end
     end
  end

endmodule
