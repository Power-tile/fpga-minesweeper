module iramHRM(CLK, RESET, ADDR, Q);
  input           CLK;
  input           RESET;
  input  [9:0]  ADDR;
  output [15:0] Q;

  reg     [15:0] mem[0:511]; // instruction memory with 16 bit entries

  wire    [8:0]  saddr;
  integer        i;


  assign saddr = ADDR[9:1];
  assign Q = mem[saddr];

  always @(posedge CLK) begin
     if(RESET) begin
        mem[0]   <= 16'b1111000000001000;    // ADD $1, $0, $0
        mem[1]   <= 16'b1111000000010000;    // ADD $2, $0, $0
        mem[2]   <= 16'b1111000000011000;    // ADD $3, $0, $0
        mem[3]   <= 16'b1001000011000001;    // BNE $3, $0, skip_jump_end[1]
        mem[4]   <= 16'b0001000010001001;    // JUMP end[137]
        mem[5]   <= 16'b0101000100000001;    // ADDI $4, $0, 1
        mem[6]   <= 16'b1111000000101000;    // ADD $5, $0, $0
        mem[7]   <= 16'b0101000111011110;    // ADDI $7, $0, 30
        mem[8]   <= 16'b0101111111011110;    // ADDI $7, $7, 30
        mem[9]   <= 16'b0101111111000100;    // ADDI $7, $7, 4
        mem[10]  <= 16'b1001111101000001;    // BNE $5, $7, skip_jump_for_end[1]
        mem[11]  <= 16'b0001000000100010;    // JUMP for_end[34]
        mem[12]  <= 16'b0101101111011110;    // ADDI $7, $5, 30
        mem[13]  <= 16'b0101111111011110;    // ADDI $7, $7, 30
        mem[14]  <= 16'b0101111111000100;    // ADDI $7, $7, 4
        mem[15]  <= 16'b0010111111000000;    // LB $7, 0($7)
        mem[16]  <= 16'b1111111000111100;    // SLL $7, $7
        mem[17]  <= 16'b1111111000111011;    // SRL $7, $7
        mem[18]  <= 16'b0101000110010000;    // ADDI $6, $0, 16
        mem[19]  <= 16'b0101110110010000;    // ADDI $6, $6, 16
        mem[20]  <= 16'b1000110111001001;    // BEQ $7, $6, first_if[9]
        mem[21]  <= 16'b0101000110011110;    // ADDI $6, $0, 30
        mem[22]  <= 16'b0101110110011110;    // ADDI $6, $6, 30
        mem[23]  <= 16'b0101110110000011;    // ADDI $6, $6, 3
        mem[24]  <= 16'b1001110111000111;    // BNE $7, $6, first_else[7]
        mem[25]  <= 16'b0010101111000000;    // LB $7, 0($5)
        mem[26]  <= 16'b0101000110011110;    // ADDI $6, $0, 30
        mem[27]  <= 16'b0101110110011110;    // ADDI $6, $6, 30
        mem[28]  <= 16'b0101110110011100;    // ADDI $6, $6, 28
        mem[29]  <= 16'b1001110111000010;    // BNE $7, $6, first_else[2]
        mem[30]  <= 16'b1111000000100000;    // ADD $4, $0, $0
        mem[31]  <= 16'b0001000000100010;    // JUMP for_end[34]
        mem[32]  <= 16'b0101101101000001;    // ADDI $5, $5, 1
        mem[33]  <= 16'b0001000000000111;    // JUMP for[7]
        mem[34]  <= 16'b1000000011000001;    // BEQ $3, $0, continue_main_if[1]
        mem[35]  <= 16'b0001000010001001;    // JUMP main_else[137]
        mem[36]  <= 16'b1001000100000001;    // BNE $4, $0, continue_mini_if[1]
        mem[37]  <= 16'b0001000000000011;    // JUMP while[3]
        mem[38]  <= 16'b1111001000111011;    // SRL $7, $1
        mem[39]  <= 16'b1111111000111011;    // SRL $7, $7
        mem[40]  <= 16'b1111111000111011;    // SRL $7, $7
        mem[41]  <= 16'b1111111000111011;    // SRL $7, $7
        mem[42]  <= 16'b1111111010111000;    // ADD $7, $7, $2
        mem[43]  <= 16'b0010111101000000;    // LB $5, 0($7)
        mem[44]  <= 16'b0101000110111111;    // ADDI $6, $0, -1
        mem[45]  <= 16'b1111110000110011;    // SRL $6, $6
        mem[46]  <= 16'b1111101110101101;    // AND $5, $5, $6
        mem[47]  <= 16'b0100111101000000;    // SB $5, 0($7)
        mem[48]  <= 16'b0101000111000111;    // ADDI $7, $0, 7
        mem[49]  <= 16'b1001111100000100;    // BNE $4, $7, elif_1[4]
        mem[50]  <= 16'b0101010111111111;    // ADDI $7, $2, -1
        mem[51]  <= 16'b1011111000000010;    // BLTZ $7, elif_1[2]
        mem[52]  <= 16'b0101010010111111;    // ADDI $2, $2, -1
        mem[53]  <= 16'b0001000001110011;    // JUMP elif_done[115]
        mem[54]  <= 16'b0101000111000101;    // ADDI $7, $0, 5
        mem[55]  <= 16'b1001111100000100;    // BNE $4, $7, elif_2[4]
        mem[56]  <= 16'b0101010111110001;    // ADDI $7, $2, -15
        mem[57]  <= 16'b1010111000000010;    // BGEZ $7, elif_2[2]
        mem[58]  <= 16'b0101010010000001;    // ADDI $2, $2, 1
        mem[59]  <= 16'b0001000001110011;    // JUMP elif_done[115]
        mem[60]  <= 16'b0101000111000100;    // ADDI $7, $0, 4
        mem[61]  <= 16'b1001111100000100;    // BNE $4, $7, elif_3[4]
        mem[62]  <= 16'b0101001111111111;    // ADDI $7, $1, -1
        mem[63]  <= 16'b1011111000000010;    // BLTZ $7, elif_3[2]
        mem[64]  <= 16'b0101001001111111;    // ADDI $1, $1, -1
        mem[65]  <= 16'b0001000001110011;    // JUMP elif_done[115]
        mem[66]  <= 16'b0101000111000110;    // ADDI $7, $0, 6
        mem[67]  <= 16'b1001111100000100;    // BNE $4, $7, elif_4[4]
        mem[68]  <= 16'b0101001111111101;    // ADDI $7, $1, -3
        mem[69]  <= 16'b1010111000000010;    // BGEZ $7, elif_4[2]
        mem[70]  <= 16'b0101001001000001;    // ADDI $1, $1, 1
        mem[71]  <= 16'b0001000001110011;    // JUMP elif_done[115]
        mem[72]  <= 16'b0101000111000001;    // ADDI $7, $0, 1
        mem[73]  <= 16'b1000111100000001;    // BEQ $4, $7, continue_elif_4[1]
        mem[74]  <= 16'b0001000001100100;    // JUMP elif_5[100]
        mem[75]  <= 16'b1111001000111011;    // SRL $7, $1
        mem[76]  <= 16'b1111111000111011;    // SRL $7, $7
        mem[77]  <= 16'b1111111000111011;    // SRL $7, $7
        mem[78]  <= 16'b1111111000111011;    // SRL $7, $7
        mem[79]  <= 16'b1111111010111000;    // ADD $7, $7, $2
        mem[80]  <= 16'b0010111110000000;    // LB $6, 0($7)
        mem[81]  <= 16'b1111110000110100;    // SLL $6, $6
        mem[82]  <= 16'b1111110000110011;    // SRL $6, $6
        mem[83]  <= 16'b0101110110100010;    // ADDI $6, $6, -30
        mem[84]  <= 16'b0101110110100010;    // ADDI $6, $6, -30
        mem[85]  <= 16'b0101110110111101;    // ADDI $6, $6, -3
        mem[86]  <= 16'b1001000110000100;    // BNE $6, $0, not_question[4]
        mem[87]  <= 16'b0101000110010000;    // ADDI $6, $0, 16
        mem[88]  <= 16'b0101110110010000;    // ADDI $6, $6, 16
        mem[89]  <= 16'b0100111110000000;    // SB $6, 0($7)
        mem[90]  <= 16'b0001000001110011;    // JUMP elif_done[115]
        mem[91]  <= 16'b0010111110000000;    // LB $6 0($7)
        mem[92]  <= 16'b0101110110110000;    // ADDI $6, $6, -16
        mem[93]  <= 16'b0101110110110000;    // ADDI $6, $6, -16
        mem[94]  <= 16'b1001000110000101;    // BNE $6, $0, elif_5[5]
        mem[95]  <= 16'b0101000110011110;    // ADDI $6, $0, 30
        mem[96]  <= 16'b0101110110011110;    // ADDI $6, $6, 30
        mem[97]  <= 16'b0101110110000011;    // ADDI $6, $6, 3
        mem[98]  <= 16'b0100111110000000;    // SB $6, 0($7)
        mem[99]  <= 16'b0001000001110011;    // JUMP elif_done[115]
        mem[100] <= 16'b0101000111000010;    // ADDI $7, $0, 2
        mem[101] <= 16'b1001111100001101;    // BNE $4, $7, elif_done[13]
        mem[102] <= 16'b1111001000111011;    // SRL $7, $1
        mem[103] <= 16'b1111111000111011;    // SRL $7, $7
        mem[104] <= 16'b1111111000111011;    // SRL $7, $7
        mem[105] <= 16'b1111111000111011;    // SRL $7, $7
        mem[106] <= 16'b1111111010111000;    // ADD $7, $7, $2
        mem[107] <= 16'b0101111111011110;    // ADDI $7, $7, 30
        mem[108] <= 16'b0101111111011110;    // ADDI $7, $7, 30
        mem[109] <= 16'b0101111111000010;    // ADDI $7, $7, 2
        mem[110] <= 16'b0010111110000000;    // LB $6 0($7)
        mem[111] <= 16'b0101111111100010;    // ADDI $7, $7, -30
        mem[112] <= 16'b0101111111100010;    // ADDI $7, $7, -30
        mem[113] <= 16'b0101111111111110;    // ADDI $7, $7, -2
        mem[114] <= 16'b0100111110000000;    // SB $6, 0($7)
        mem[115] <= 16'b1111001000111011;    // SRL $7, $1
        mem[116] <= 16'b1111111000111011;    // SRL $7, $7
        mem[117] <= 16'b1111111000111011;    // SRL $7, $7
        mem[118] <= 16'b1111111000111011;    // SRL $7, $7
        mem[119] <= 16'b1111111010111000;    // ADD $7, $7, $2
        mem[120] <= 16'b0010111110000000;    // LB $6, 0($7)
        mem[121] <= 16'b0111110110111111;    // ORI $6, $6, -1
        mem[122] <= 16'b0100111110000000;    // SB $6, 0($7)
        mem[123] <= 16'b1111001000111011;    // SRL $7, $1
        mem[124] <= 16'b1111111000111011;    // SRL $7, $7
        mem[125] <= 16'b1111111000111011;    // SRL $7, $7
        mem[126] <= 16'b1111111000111011;    // SRL $7, $7
        mem[127] <= 16'b1111111010111000;    // ADD $7, $7, $2
        mem[128] <= 16'b1111110000110100;    // SLL $6, $6
        mem[129] <= 16'b1111110000110011;    // SRL $6, $6
        mem[130] <= 16'b0010111110000000;    // LB $6, 0($7)
        mem[131] <= 16'b0101000111011110;    // ADDI $7, $0, 30
        mem[132] <= 16'b0101000111011110;    // ADDI $7, $0, 30
        mem[133] <= 16'b0101000111011100;    // ADDI $7, $0, 28
        mem[134] <= 16'b1001111110000001;    // BNE $6, $7, not_dead[1]
        mem[135] <= 16'b0101000011000001;    // ADDI $3, $0, 1
        mem[136] <= 16'b0001000000000011;    // JUMP while[3]
        mem[137] <= 16'b0000000000000001;    // HALT

        for(i = 138; i < 512; i = i + 1) begin
          mem[i] <= 16'b0000000000000000;
        end
     end
  end

endmodule
